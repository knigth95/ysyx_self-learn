module top(
    init begin:
        $display("Hello, world!");
        $finish;
    end
    );
endmodule
