module top(a,b,f);
  input [3:0]a;
endmodule