module top(;
    initial begin:
        $display("Hello, world!");
        $finish;
    end
    );
endmodule
