module example(
   input a,
   input b,
   input f
);
     
     
  endmodule
