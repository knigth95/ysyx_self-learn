module example(
   input a,
   input;
);
     
     
  endmodule
