module example;
     
     
  endmodule
