module top:
    