module example(
   input a,
   ;
);
     
     
  endmodule
