module example(
   input a,
   input b,
   put f
);
   assign f=a^b;
endmodule
