module top(
     begin:
        $display("Hello, world!");
        $finish;
    end
    );
endmodule
