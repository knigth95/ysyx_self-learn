module top(a,b,f);

endmodule