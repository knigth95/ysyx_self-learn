module top:
    initial begin:
    