module top:
