module example(
   input a,
   input b;
);
     
     
  endmodule
