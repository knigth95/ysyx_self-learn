module example(
   input ;
);
     
     
  endmodule
