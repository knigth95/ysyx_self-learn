module top(a,b,f);
  
  assi
endmodule