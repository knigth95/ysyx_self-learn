module example(
   
);
     
     
  endmodule
