module top(a,b,f);
  input [];
endmodule