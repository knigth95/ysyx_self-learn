module example(
   input a,
   input b,
   input f
);
   assign f=a^b;
endmodule
