module ex;
     initial begin $display("Hello World"); $finish; end
  endmodule
