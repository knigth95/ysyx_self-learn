module top(
    in begin:
        $display("Hello, world!");
        $finish;
    end
    );
endmodule
