module top(a,b,c);

endmodule