module top(a,);

endmodule