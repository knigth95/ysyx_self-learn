module example;
     
     end
  endmodule
